package rutr_pkg;

import uvm_pkg::*;

`include "uvm_macros.svh"

`include "source_agt_config.sv"
`include "dest_agt_config.sv"
`include "rutr_env_config.sv"

`include "source_xtn.sv"
`include "source_driver.sv"
`include "source_sequencer.sv"
`include "source_monitor.sv"
`include "source_agt.sv"
`include "source_agt_top.sv"
`include "source_sequence.sv"

`include "dest_xtn.sv"
`include "dest_driver.sv"
`include "dest_monitor.sv"
`include "dest_sequencer.sv"
`include "dest_agt.sv"
`include "dest_agt_top.sv"
`include "dest_sequence.sv"

`include " rutr_scoreboard.sv"

`include "rutr_env.sv"
`include "rutr_test.sv"


endpackage

